library verilog;
use verilog.vl_types.all;
entity mic1 is
    port(
        \00\            : out    vl_logic;
        \10\            : in     vl_logic;
        \11\            : in     vl_logic;
        \01\            : out    vl_logic;
        \02\            : out    vl_logic;
        \03\            : out    vl_logic
    );
end mic1;
